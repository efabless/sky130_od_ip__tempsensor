** sch_path: /home/tim/gits/chipalooza_projects_redef/dependencies/sky130_od_ip__tempsensor/xschem/sky130_od_ip__tempsensor_ext_vp.sch
.subckt sky130_od_ip__tempsensor_ext_vp vbe1_out vdd vss vbg ena vbe2_out
*.PININFO vdd:I vss:I vbe2_out:O vbe1_out:O ena:I vbg:I
XQ_BL1 vss vss vbe1 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ_BR1 vss vss vbe2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XM4 net2 vbg net1 vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM5 vp vp net1 vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM7 vp net2 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM8 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM3 vp ena vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 m=1
XM6 net1 ena vss vss sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
x1 vdd vss ena vbe1 vbe1_out buffer
x2 vdd vss ena vbe2 vbe2_out buffer
XM1 vbe1 vp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=1
XM2 vbe2 vp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 m=5
XD1 vss ena sky130_fd_pr__diode_pw2nd_05v5 area=202.5e11 perim=1.8e6
XD2 vss vbg sky130_fd_pr__diode_pw2nd_05v5 area=202.5e11 perim=1.8e6
XD3 vss vbe1 sky130_fd_pr__diode_pw2nd_05v5 area=202.5e11 perim=1.8e6
XD4 vss vbe2 sky130_fd_pr__diode_pw2nd_05v5 area=202.5e11 perim=1.8e6
.ends

* expanding   symbol:  buffer.sym # of pins=5
** sym_path: /home/tim/gits/chipalooza_projects_redef/dependencies/sky130_od_ip__tempsensor/xschem/buffer.sym
** sch_path: /home/tim/gits/chipalooza_projects_redef/dependencies/sky130_od_ip__tempsensor/xschem/buffer.sch
.subckt buffer vdd vss vbias input output
*.PININFO output:O input:I vdd:I vss:I vbias:I
XM1 net2 input net1 vss sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
XM2 output output net1 vss sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
XM5 net1 vbias vss vss sky130_fd_pr__nfet_01v8 L=10 W=1 nf=1 m=1
XM4 output net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=10 W=1 nf=1 m=1
XM3 net2 net2 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=10 W=1 nf=1 m=1
.ends

.end
