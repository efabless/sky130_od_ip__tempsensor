** sch_path: /home/azwefabless/cheetah_v3_analog/dependencies/sky130_od_ip__tempsensor/xschem/sky130_od_ip__tempsensor.sch
.subckt sky130_od_ip__tempsensor vdd vss Vbe2 Vbe1 ena
*.PININFO vdd:I vss:I Vbe2:O Vbe1:O ena:I
XM12 net1 Vp vdd vdd sky130_fd_pr__pfet_01v8 L=5.0 W=1 nf=1 m=5
XM13 net2 Vp vdd vdd sky130_fd_pr__pfet_01v8 L=5.0 W=1 nf=1 m=1
XQ_BR vss net10 net1 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ_BL vss vss net3 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XM11 net4 Vp vdd vdd sky130_fd_pr__pfet_01v8 L=5.0 W=1 nf=1 m=2
XM6 net5 net2 net4 net4 sky130_fd_pr__pfet_01v8 L=5.0 W=1 nf=1 m=1
XM5 net6 net1 net4 net4 sky130_fd_pr__pfet_01v8 L=5.0 W=1 nf=1 m=1
XM2 net5 net5 vss vss sky130_fd_pr__nfet_01v8 L=10.0 W=1 nf=1 m=1
XM1 net6 net6 vss vss sky130_fd_pr__nfet_01v8 L=10.0 W=1 nf=1 m=1
XM9 net7 Vp vdd vdd sky130_fd_pr__pfet_01v8 L=5.0 W=1 nf=1 m=1
XM10 Vp Vp vdd vdd sky130_fd_pr__pfet_01v8 L=5.0 W=1 nf=1 m=4
XM7 Vp net7 net9 net9 sky130_fd_pr__nfet_01v8 L=5.0 W=1 nf=1 m=4
XM8 net7 net7 net8 net8 sky130_fd_pr__nfet_01v8 L=5.0 W=1 nf=1 m=1
XM3 net9 net5 vss vss sky130_fd_pr__nfet_01v8 L=10.0 W=1 nf=1 m=4
XM4 net8 net8 vss vss sky130_fd_pr__nfet_01v8 L=5.0 W=1 nf=1 m=1
XQ_BL1 vss vss Vbe1 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ_BR1 vss vss Vbe2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XM14 Vbe1 Vp vdd vdd sky130_fd_pr__pfet_01v8 L=5.0 W=1 nf=1 m=1
XM15 Vbe2 Vp vdd vdd sky130_fd_pr__pfet_01v8 L=5.0 W=1 nf=1 m=5
XM16 Vp ena vdd vdd sky130_fd_pr__pfet_01v8 L=1.2 W=10 nf=1 m=1
R1 net3 net2 sky130_fd_pr__res_generic_l1 W=1 L=1000 m=1
R2 vss net10 sky130_fd_pr__res_generic_l1 W=1 L=200 m=1
.ends
.end
