magic
tech sky130A
magscale 1 2
timestamp 1713290077
<< pwell >>
rect 2316 -1858 4154 -1856
rect 2006 -1954 4154 -1858
<< locali >>
rect 746 432 5440 496
rect 746 328 1134 432
rect 5338 328 5440 432
rect 746 180 5440 328
rect 3018 -816 3122 -596
rect 3018 -848 3124 -816
rect 3020 -1106 3124 -848
rect 3014 -1108 3124 -1106
rect 3006 -1110 3124 -1108
rect 4264 -1110 5412 -1108
rect 726 -1304 5412 -1110
rect 726 -1470 1020 -1304
rect 1870 -1410 5412 -1304
rect 1870 -1470 2018 -1410
rect 726 -1532 2018 -1470
rect 726 -1710 2126 -1532
rect 4254 -1708 5412 -1410
rect 726 -1760 2018 -1710
rect 726 -1858 2014 -1760
rect 4264 -1852 5412 -1708
rect 4012 -1856 5412 -1852
rect 2316 -1858 5412 -1856
rect 726 -1938 5412 -1858
rect 726 -1950 4338 -1938
rect 726 -1954 4154 -1950
rect 726 -1956 812 -1954
<< viali >>
rect 1134 328 5338 432
rect 1020 -1470 1870 -1304
<< metal1 >>
rect 810 470 1092 476
rect 810 432 5400 470
rect 810 328 1134 432
rect 5338 328 5400 432
rect 810 294 5400 328
rect 810 266 1092 294
rect 1142 44 2786 124
rect 778 42 2786 44
rect 774 -136 2786 42
rect 3038 34 3158 294
rect 774 -142 940 -136
rect 774 -806 842 -142
rect 1142 -236 2786 -136
rect 2966 -142 3228 34
rect 3514 -232 4954 124
rect 5254 -142 5430 36
rect 2506 -304 2780 -236
rect 3518 -304 3704 -232
rect 1138 -580 1338 -380
rect 2502 -498 3706 -304
rect 5134 -372 5256 -370
rect 5292 -372 5426 -142
rect 2506 -500 2780 -498
rect 5134 -572 5430 -372
rect 1142 -728 1336 -580
rect 772 -974 916 -806
rect 774 -976 842 -974
rect 1138 -1064 2640 -728
rect 3464 -806 4966 -728
rect 5134 -806 5256 -572
rect 3018 -810 3120 -808
rect 2942 -986 3202 -810
rect 3018 -1198 3120 -986
rect 3464 -992 5262 -806
rect 3464 -1064 4966 -992
rect 754 -1246 1890 -1244
rect 754 -1304 1912 -1246
rect 754 -1334 1020 -1304
rect 752 -1402 1020 -1334
rect 754 -1470 1020 -1402
rect 1870 -1470 1912 -1304
rect 3018 -1332 4374 -1198
rect 754 -1536 1912 -1470
rect 754 -1538 1890 -1536
rect 756 -1772 1898 -1582
rect 2402 -1772 3814 -1454
rect 4268 -1532 4374 -1332
rect 4154 -1710 4374 -1532
rect 756 -1852 3816 -1772
rect 756 -1856 1898 -1852
use sky130_fd_pr__nfet_01v8_QXBCRM  XM1 paramcells
timestamp 1713290077
transform 1 0 1929 0 1 -898
box -1196 -310 1196 310
use sky130_fd_pr__nfet_01v8_QXBCRM  XM2
timestamp 1713290077
transform 1 0 4215 0 1 -898
box -1196 -310 1196 310
use sky130_fd_pr__pfet_01v8_lvt_B5H3CA  XM3 paramcells
timestamp 1713290077
transform 1 0 1955 0 1 -55
box -1196 -319 1196 319
use sky130_fd_pr__pfet_01v8_lvt_B5H3CA  XM4
timestamp 1713290077
transform 1 0 4241 0 1 -55
box -1196 -319 1196 319
use sky130_fd_pr__nfet_01v8_QXBCRM  XM5
timestamp 1713290077
transform 1 0 3141 0 1 -1622
box -1196 -310 1196 310
<< labels >>
flabel metal1 792 -1470 992 -1270 0 FreeSans 256 0 0 0 vss
port 1 nsew
flabel metal1 818 268 1018 468 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 5230 -572 5430 -372 0 FreeSans 256 0 0 0 output
port 4 nsew
flabel metal1 1138 -580 1338 -380 0 FreeSans 256 0 0 0 input
port 3 nsew
flabel metal1 792 -1798 992 -1598 0 FreeSans 256 0 0 0 vbias
port 2 nsew
<< end >>
