* NGSPICE file created from sky130_od_ip__tempsensor_ext_vp.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_QXBCRM a_n1000_n188# a_n1160_n274# a_1000_n100# a_n1058_n100#
X0 a_1000_n100# a_n1000_n188# a_n1058_n100# a_n1160_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_B5H3CA w_n1196_n319# a_n1000_n197# a_1000_n100#
+ a_n1058_n100#
X0 a_1000_n100# a_n1000_n197# a_n1058_n100# w_n1196_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=10
.ends

.subckt buffer input output vbias vss vdd
XXM1 input vss m1_2942_n986# m1_772_n974# sky130_fd_pr__nfet_01v8_QXBCRM
XXM2 output vss output m1_2942_n986# sky130_fd_pr__nfet_01v8_QXBCRM
XXM3 vdd m1_772_n974# vdd m1_772_n974# sky130_fd_pr__pfet_01v8_lvt_B5H3CA
XXM4 vdd m1_772_n974# output vdd sky130_fd_pr__pfet_01v8_lvt_B5H3CA
XXM5 vbias vss m1_2942_n986# vss sky130_fd_pr__nfet_01v8_QXBCRM
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_FT76RJ a_n147_n147# a_n45_n45#
X0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 perim=1.8e+06 area=2.025e+11
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_6VRZAW a_100_n536# w_n296_n1191# a_n100_675# a_100_336#
+ a_n158_n536# a_n158_772# a_n100_n633# a_n100_239# a_n100_n197# a_100_n100# a_n158_336#
+ a_100_n972# a_n158_n100# a_100_772# a_n158_n972# a_n100_n1069#
X0 a_100_336# a_n100_239# a_n158_336# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X1 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X2 a_100_772# a_n100_675# a_n158_772# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X3 a_100_n536# a_n100_n633# a_n158_n536# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
X4 a_100_n972# a_n100_n1069# a_n158_n972# w_n296_n1191# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_3VR9VM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_3HMWVM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_69TQ3K a_n260_n274# a_100_n100# a_n158_n100# a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n260_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_od_ip__tempsensor_ext_vp vdd vss vbe2_out vbe1_out ena vbg
Xx1 x1/input vbe2_out ena vss vdd buffer
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_1 vss ena sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0 vss vbg sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xx2 x2/input vbe1_out ena vss vdd buffer
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_2 vss vbe1_out sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
Xsky130_fd_pr__diode_pw2nd_05v5_FT76RJ_3 vss vbe2_out sky130_fd_pr__diode_pw2nd_05v5_FT76RJ
XXQ_BR1 x1/input vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXQ_BL1 x2/input vss vss sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
XXM22 vdd vdd vp vdd x1/input x1/input vp vp vp vdd x1/input vdd x1/input vdd x1/input
+ vp sky130_fd_pr__pfet_01v8_lvt_6VRZAW
XXM11 vdd vp vdd x2/input sky130_fd_pr__pfet_01v8_lvt_3VR9VM
XXM33 vdd ena vp vdd sky130_fd_pr__pfet_01v8_3HMWVM
XXM44 vss m1_772_n1144# m1_420_n380# vbg sky130_fd_pr__nfet_01v8_69TQ3K
XXM55 vss vp m1_772_n1144# vp sky130_fd_pr__nfet_01v8_69TQ3K
XXM66 ena vss m1_772_n1144# vss sky130_fd_pr__nfet_01v8_QXBCRM
XXM77 vdd m1_420_n380# vp vdd sky130_fd_pr__pfet_01v8_3HMWVM
XXM88 vdd m1_420_n380# vdd m1_420_n380# sky130_fd_pr__pfet_01v8_3HMWVM
.ends

